//-----------------------------------------------------------------
module SHIFTER_RIGHT_16BITS (in, s, out);
    input wire [15:0] in;
    input wire [3:0] s;
    output wire [15:0] out;
    wire [15:0] net0, net1, net2;

//--1BIT-----------------------------------------------------
mux2X16 entity_1 (in, {1'b0,in[15:1]}, s[0], net0);
//--2BITS----------------------------------------------------
mux2X16 entity_2 (net0, {2'b0,net0[15:2]}, s[1], net1);
//--4BITS---------------------------------------------------
mux2X16 entity_3 (net1, {4'b0,net1[15:4]}, s[2], net2);
//--8BITS---------------------------------------------------
mux2X16 entity_4 (net2, {8'b0,net2[15:8]}, s[3], out);
endmodule
//-----------------------------------------------------------------
module SHIFTER_RIGHT_24BITS (in, s, out);
    input wire [23:0] in;
    input wire [4:0] s;
    output wire [23:0] out;
    wire [23:0] net0, net1, net2, net3;

//--1BIT-----------------------------------------------------
mux2X24 entity_5 (in, {1'b0,in[23:1]}, s[0], net0);
//--2BITS----------------------------------------------------
mux2X24 entity_6 (net0, {2'b0,net0[23:2]}, s[1], net1);
//--4BITS---------------------------------------------------
mux2X24 entity_7 (net1, {4'b0,net1[23:4]}, s[2], net2);
//--8BITS---------------------------------------------------
mux2X24 entity_8 (net2, {8'b0,net2[23:8]}, s[3], net3);
//--16BITS-------------------------------------------------
mux2X24 entity_9 (net3, {16'b0,net3[23:16]}, s[4], out);
endmodule
//-----------------------------------------------------------------
module SHIFTER_RIGHT_32BITS (in, s, out);

    input wire [31:0] in;
    input wire [4:0] s;
    output wire [31:0] out;
    wire [31:0] net0, net1, net2, net3;

//--1BIT-----------------------------------------------------
mux2X32 entity_10 (in, {1'b0,in[31:1]}, s[0], net0);
//--2BITS----------------------------------------------------
mux2X32 entity_11 (net0, {2'b0,net0[31:2]}, s[1], net1);
//--4BITS---------------------------------------------------
mux2X32 entity_12 (net1, {4'b0,net1[31:4]}, s[2], net2);
//--8BITS---------------------------------------------------
mux2X32 entity_13 (net2, {8'b0,net2[31:8]}, s[3], net3);
//--16BITS-------------------------------------------------
mux2X32 entity_14 (net3, {16'b0,net3[31:16]}, s[4], out);
endmodule
//----------------------------------------------------------
module SHIFTER_RIGHT_48BITS (in, s, out);
    input wire [47:0] in;
    input wire [5:0] s;
    output wire [47:0] out;
    wire [47:0] net0, net1, net2, net3, net4;
//--1BIT-----------------------------------------------------
mux2X48 entity_15 (in, {1'b0,in[47:1]}, s[0], net0);
//--2BITS----------------------------------------------------
mux2X48 entity_16 (net0, {2'b0,net0[47:2]}, s[1], net1);
//--4BITS---------------------------------------------------
mux2X48 entity_17 (net1, {4'b0,net1[47:4]}, s[2], net2);
//--8BITS---------------------------------------------------
mux2X48 entity_18 (net2, {8'b0,net2[47:8]}, s[3], net3);
//--16BITS-------------------------------------------------
mux2X48 entity_19 (net3, {16'b0,net3[47:16]}, s[4], net4);
//--32BITS-------------------------------------------------
mux2X48 entity_10 (net4, {32'b0,net4[47:32]}, s[5], out);
endmodule
//----------------------------------------------------------
module SHIFTER_RIGHT_64BITS (in, s, out);
    input wire [63:0] in;
    input wire [5:0] s;
    output wire [63:0] out;
    wire [63:0] net0, net1, net2, net3, net4;
//--1BIT-----------------------------------------------------
mux2X64 entity_11 (in, {1'b0,in[63:1]}, s[0], net0);
//--2BITS----------------------------------------------------
mux2X64 entity_12 (net0, {2'b0,net0[63:2]}, s[1], net1);
//--4BITS---------------------------------------------------
mux2X64 entity_13 (net1, {4'b0,net1[63:4]}, s[2], net2);
//--8BITS---------------------------------------------------
mux2X64 entity_14 (net2, {8'b0,net2[63:8]}, s[3], net3);
//--16BITS-------------------------------------------------
mux2X64 entity_15 (net3, {16'b0,net3[63:16]}, s[4], net4);
//--32BITS-------------------------------------------------
mux2X64 entity_16 (net4, {32'b0,net4[63:32]}, s[5], out);
endmodule
//----------------------------------------------------------

`timescale 1ns/1ps
module SHIFTER_RIGHT_BITS_TB;
    reg [47:0] a;
    reg [5:0] b;
    wire [47:0] c;

SHIFTER_RIGHT_48BITS uut (a, b, c);
    initial begin
        #10
        a = 48'd10000000;
        b = 6'd10;
        #10
        a = 48'd65400000;
        b = 6'd9;
        #10
        a = 48'd1230124;
        b = 6'd3;

    end
endmodule
