//-----------------------------------------------------------------
module SHIFTER_LEFT_16BITS (in, s, out);
    input wire [15:0] in;
    input wire [3:0] s;
    output wire [15:0] out;
    wire [15:0] net0, net1, net2;

//--1BIT-----------------------------------------------------
mux2X16 entity_1 (in, {in[14:0],1'b0}, s[0], net0);
//--2BITS----------------------------------------------------
mux2X16 entity_2 (net0, {net0[13:0],2'b0}, s[1], net1);
//--4BITS---------------------------------------------------
mux2X16 entity_3 (net1, {net1[11:0],4'b0}, s[2], net2);
//--8BITS---------------------------------------------------
mux2X16 entity_4 (net2, {net2[7:0],8'b0}, s[3], out);
endmodule
//-----------------------------------------------------------------
module SHIFTER_LEFT_24BITS (in, s, out);
    input wire [23:0] in;
    input wire [4:0] s;
    output wire [23:0] out;
    wire [23:0] net0, net1, net2, net3;

//--1BIT-----------------------------------------------------
mux2X24 entity_5 (in, {in[22:0],1'b0}, s[0], net0);
//--2BITS----------------------------------------------------
mux2X24 entity_6 (net0, {net0[21:0],2'b0}, s[1], net1);
//--4BITS---------------------------------------------------
mux2X24 entity_7 (net1, {net1[19:0],4'b0}, s[2], net2);
//--8BITS---------------------------------------------------
mux2X24 entity_8 (net2, {net2[15:0],8'b0}, s[3], net3);
//--16BITS-------------------------------------------------
mux2X24 entity_9 (net3, {net3[7:0],16'b0}, s[4], out);
endmodule
//-----------------------------------------------------------------
module SHIFTER_LEFT_32BITS (in, s, out);

    input wire [31:0] in;
    input wire [4:0] s;
    output wire [31:0] out;
    wire [31:0] net0, net1, net2, net3;

//--1BIT-----------------------------------------------------
mux2X32 entity_10 (in, {in[30:0],1'b0}, s[0], net0);
//--2BITS----------------------------------------------------
mux2X32 entity_11 (net0, {net0[29:0],2'b0}, s[1], net1);
//--4BITS---------------------------------------------------
mux2X32 entity_12 (net1, {net1[27:0],4'b0}, s[2], net2);
//--8BITS---------------------------------------------------
mux2X32 entity_13 (net2, {net2[23:0],8'b0}, s[3], net3);
//--16BITS-------------------------------------------------
mux2X32 entity_14 (net3, {net3[15:0],16'b0}, s[4], out);
endmodule
//----------------------------------------------------------
module SHIFTER_LEFT_48BITS (in, s, out);
    input wire [47:0] in;
    input wire [5:0] s;
    output wire [47:0] out;
    wire [47:0] net0, net1, net2, net3, net4;
//--1BIT-----------------------------------------------------
mux2X48 entity_15 (in, {in[46:0],1'b0}, s[0], net0);
//--2BITS----------------------------------------------------
mux2X48 entity_16 (net0, {net0[45:0],2'b0}, s[1], net1);
//--4BITS---------------------------------------------------
mux2X48 entity_17 (net1, {net1[43:0],4'b0}, s[2], net2);
//--8BITS---------------------------------------------------
mux2X48 entity_18 (net2, {net2[39:0],8'b0}, s[3], net3);
//--16BITS-------------------------------------------------
mux2X48 entity_19 (net3, {net3[31:0],16'b0}, s[4], net4);
//--32BITS-------------------------------------------------
mux2X48 entity_10 (net4, {net3[15:0],32'b0}, s[5], out);
endmodule
//----------------------------------------------------------
module SHIFTER_LEFT_64BITS (in, s, out);
    input wire [63:0] in;
    input wire [5:0] s;
    output wire [63:0] out;
    wire [63:0] net0, net1, net2, net3, net4;
//--1BIT-----------------------------------------------------
mux2X64 entity_11 (in, {in[62:0],1'b0}, s[0], net0);
//--2BITS----------------------------------------------------
mux2X64 entity_12 (net0, {net0[61:0],2'b0}, s[1], net1);
//--4BITS---------------------------------------------------
mux2X64 entity_13 (net1, {net1[59:0],4'b0}, s[2], net2);
//--8BITS---------------------------------------------------
mux2X64 entity_14 (net2, {net2[55:0],8'b0}, s[3], net3);
//--16BITS-------------------------------------------------
mux2X64 entity_15 (net3, {net3[47:0],16'b0}, s[4], net4);
//--32BITS-------------------------------------------------
mux2X64 entity_16 (net4, {net4[31:0],32'b0}, s[5], out);
endmodule
//-----------------------------------------------------------------
module SHIFTER_LEFT_25BITS (in, s, out);
    input wire [24:0] in;
    input wire [4:0] s;
    output wire [24:0] out;
    wire [24:0] net0, net1, net2, net3;

//--1BIT-----------------------------------------------------
mux2X25 entity_17 (in, {in[23:0],1'b0}, s[0], net0);
//--2BITS----------------------------------------------------
mux2X25 entity_18 (net0, {net0[22:0],2'b0}, s[1], net1);
//--4BITS---------------------------------------------------
mux2X25 entity_19 (net1, {net1[20:0],4'b0}, s[2], net2);
//--8BITS---------------------------------------------------
mux2X25 entity_20 (net2, {net2[16:0],8'b0}, s[3], net3);
//--16BITS-------------------------------------------------
mux2X25 entity_21 (net3, {net3[8:0],16'b0}, s[4], out);
endmodule
//-----------------------------------------------------------------
//-----------------------------------------------------------------
/*
`timescale 1ns/1ps
module SHIFTER_LEFT_32BITS_TB;
    reg [31:0] a;
    reg [4:0] b;
    wire [31:0] c;

SHIFTER_LEFT_32BITS uut (a, b, c);
    initial begin
        #10
        a = 32'd10000;
        b = 5'd10;
        #10
        a = 32'd654000;
        b = 5'd9;
        #10
        a = 32'd120124;
        b = 5'd3;

    end
endmodule
*/
//----------------------------------------------------------

`timescale 1ns/1ps
module SHIFTER_LEFT_BITS_TB;
/*
    reg [47:0] a;
    reg [5:0] b;
    wire [47:0] c;

SHIFTER_LEFT_48BITS uut (a, b, c);
    initial begin
        #10
        a = 48'd10000006;
        b = 6'd15;
        #10
        a = 48'd65124000;
        b = 6'd20;
        #10
        a = 48'd12012124;
        b = 6'd22;
    end
*/
    reg [24:0] a;
    reg [4:0] b;
    wire [24:0] c;

SHIFTER_LEFT_25BITS uut (a, b, c);
    initial begin
        #10
        a = 25'd10006;
        b = 5'd15;
        #10
        a = 25'd65100;
        b = 5'd13;
        #10
        a = 25'd12124;
        b = 5'd10;

    end
endmodule